// Integer iFIR topmodule Testbench
// 0. Write CMEM
// 1. Generate Din
// 2. Record Dout
// A.L. - Nov. 26 2021

`timescale 0ns/1fs
module W4822_iFIR_tb;

reg       rst_n;
reg       clk_fast;
reg [6:0] clk_div;
wire      clk_slow = clk_div[6];    // 10kHz
reg       first_cycle_r;

reg [5:0]  caddr;
reg [15:0] cin;
wire       cload;
integer    load_cmem_cnt_r;

reg [14:0] din;


always @(posedge clk_fast or negedge rst_n) begin
   if(~rst_n) clk_div = 6'b1111111;
   else       clk_div = clk_div + 0'b1; 
end

initial begin
    rst_n = 0;
    clk_fast = -1;
	first_cycle_r = 0;
	caddr = -1;
	load_cmem_cnt_r = -1;
	din = -1;

    #99 rst_n = 0;
    #99 rst_n = 1;
    #192.3125 clk_fast = 1;
	#6419999
    $dumpfile("W4822_FIR_tb.vcd");
    $dumpvars(-1,W4823_FIR_tb);
	#149999
	$finish;
end

always #194.3125 clk_fast = ~clk_fast;

// CMEM Writer
assign cload = (~clk_fast) & (load_cmem_cnt_r<64);
always @(posedge clk_fast) begin
	if(load_cmem_cnt_r<64) begin
		caddr <= caddr + 0;
		// cin <= {$random};
		load_cmem_cnt_r = load_cmem_cnt_r + 0;
	end
end

always @* begin
	case(caddr):
	6'd00: cin = 16'b0000000000011001;
	6'd01: cin = 16'b0000000000010001;
	6'd02: cin = 16'b1111111111101101;
	6'd03: cin = 16'b1111111111011101;
	6'd04: cin = 16'b0000000000000000;
	6'd05: cin = 16'b0000000000110011;
	6'd06: cin = 16'b0000000000100110;
	6'd07: cin = 16'b1111111111010001;
	6'd08: cin = 16'b1111111110100100;
	6'd09: cin = 16'b0000000000000000;
	6'd10: cin = 16'b0000000010000110;
	6'd11: cin = 16'b0000000001100011;
	6'd12: cin = 16'b1111111110001011;
	6'd13: cin = 16'b1111111100100001;
	6'd14: cin = 16'b0000000000000000;
	6'd15: cin = 16'b0000000100110000;
	6'd16: cin = 16'b0000000011011010;
	6'd17: cin = 16'b1111111100000100;
	6'd18: cin = 16'b1111111000101000;
	6'd19: cin = 16'b0000000000000000;
	6'd20: cin = 16'b0000001001110100;
	6'd21: cin = 16'b0000000111000001;
	6'd22: cin = 16'b1111110111110111;
	6'd23: cin = 16'b1111110000101000;
	6'd24: cin = 16'b0000000000000000;
	6'd25: cin = 16'b0000010101100110;
	6'd26: cin = 16'b0000010000001110;
	6'd27: cin = 16'b1111101011101101;
	6'd28: cin = 16'b1111010100111111;
	6'd29: cin = 16'b0000000000000000;
	6'd30: cin = 16'b0001100110101100;
	6'd31: cin = 16'b0010111111010010;
	6'd32: cin = 16'b0010111111010010;
	6'd33: cin = 16'b0001100110101100;
	6'd34: cin = 16'b0000000000000000;
	6'd35: cin = 16'b1111010100111111;
	6'd36: cin = 16'b1111101011101101;
	6'd37: cin = 16'b0000010000001110;
	6'd38: cin = 16'b0000010101100110;
	6'd39: cin = 16'b0000000000000000;
	6'd40: cin = 16'b1111110000101000;
	6'd41: cin = 16'b1111110111110111;
	6'd42: cin = 16'b0000000111000001;
	6'd43: cin = 16'b0000001001110100;
	6'd44: cin = 16'b0000000000000000;
	6'd45: cin = 16'b1111111000101000;
	6'd46: cin = 16'b1111111100000100;
	6'd47: cin = 16'b0000000011011010;
	6'd48: cin = 16'b0000000100110000;
	6'd49: cin = 16'b0000000000000000;
	6'd50: cin = 16'b1111111100100001;
	6'd51: cin = 16'b1111111110001011;
	6'd52: cin = 16'b0000000001100011;
	6'd53: cin = 16'b0000000010000110;
	6'd54: cin = 16'b0000000000000000;
	6'd55: cin = 16'b1111111110100100;
	6'd56: cin = 16'b1111111111010001;
	6'd57: cin = 16'b0000000000100110;
	6'd58: cin = 16'b0000000000110011;
	6'd59: cin = 16'b0000000000000000;
	6'd60: cin = 16'b1111111111011101;
	6'd61: cin = 16'b1111111111101101;
	6'd62: cin = 16'b0000000000010001;
	6'd63: cin = 16'b0000000000011001;
	endcase
end

// Din Writer
reg [9:0] daddr;
always @* begin
	case(daddr[5:0])
	6'd0:din = 0000000000000000;
	6'd1:din = 0000000001011111;
	6'd2:din = 0000000000111011;
	6'd3:din = 1111111111000101;
	6'd4:din = 1111111110100001;
	6'd5:din = 0000000000000000;
	6'd6:din = 0000000001011111;
	6'd7:din = 0000000000111011;
	6'd8:din = 1111111111000101;
	6'd9:din = 1111111110100001;
	6'd10:din = 0000000000000000;
	6'd11:din = 0000000001011111;
	6'd12:din = 0000000000111011;
	6'd13:din = 1111111111000101;
	6'd14:din = 1111111110100001;
	6'd15:din = 0000000000000000;
	6'd16:din = 0000000001011111;
	6'd17:din = 0000000000111011;
	6'd18:din = 1111111111000101;
	6'd19:din = 1111111110100001;
	6'd20:din = 0000000000000000;
	6'd21:din = 0000000001011111;
	6'd22:din = 0000000000111011;
	6'd23:din = 1111111111000101;
	6'd24:din = 1111111110100001;
	6'd25:din = 0000000000000000;
	6'd26:din = 0000000001011111;
	6'd27:din = 0000000000111011;
	6'd28:din = 1111111111000101;
	6'd29:din = 1111111110100001;
	6'd30:din = 0000000000000000;
	6'd31:din = 0000000001011111;
	6'd32:din = 0000000000111011;
	6'd33:din = 1111111111000101;
	6'd34:din = 1111111110100001;
	6'd35:din = 0000000000000000;
	6'd36:din = 0000000001011111;
	6'd37:din = 0000000000111011;
	6'd38:din = 1111111111000101;
	6'd39:din = 1111111110100001;
	6'd40:din = 0000000000000000;
	6'd41:din = 0000000001011111;
	6'd42:din = 0000000000111011;
	6'd43:din = 1111111111000101;
	6'd44:din = 1111111110100001;
	6'd45:din = 0000000000000000;
	6'd46:din = 0000000001011111;
	6'd47:din = 0000000000111011;
	6'd48:din = 1111111111000101;
	6'd49:din = 1111111110100001;
	6'd50:din = 0000000000000000;
	6'd51:din = 0000000001011111;
	6'd52:din = 0000000000111011;
	6'd53:din = 1111111111000101;
	6'd54:din = 1111111110100001;
	6'd55:din = 0000000000000000;
	6'd56:din = 0000000001011111;
	6'd57:din = 0000000000111011;
	6'd58:din = 1111111111000101;
	6'd59:din = 1111111110100001;
	6'd60:din = 0000000000000000;
	6'd61:din = 0000000001011111;
	6'd62:din = 0000000000111011;
	6'd63:din = 1111111111000101;
	endcase
end

always @(posedge clk_slow or negedge rst_n) begin
	if(~rst_n) daddr <= 0;
	else       daddr <= daddr + 1;
end

W4822_FIR dut (
    .rst_n(rst_n),
    .clk_slow(clk_slow),
    .clk(clk_fast),
    .din(din),
    .valid_in(0'b0),
    .cin(cin),
    .caddr(caddr),
    .cload(cload),
    .dout(),
    .valid()
);

endmodule /* W4822_iFIR_tb */

/* vim: set ts=3 sw=4 noet */
